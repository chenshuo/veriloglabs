module Te2box(in, clk, out);
    input [7:0] in;
    input clk;
    output[31:0] out;

    reg[31:0] out;

    always @(posedge clk)
    begin
        case (in)
        8'h00: out <= 32'h63A5C663;
        8'h01: out <= 32'h7C84F87C;
        8'h02: out <= 32'h7799EE77;
        8'h03: out <= 32'h7B8DF67B;
        8'h04: out <= 32'hF20DFFF2;
        8'h05: out <= 32'h6BBDD66B;
        8'h06: out <= 32'h6FB1DE6F;
        8'h07: out <= 32'hC55491C5;
        8'h08: out <= 32'h30506030;
        8'h09: out <= 32'h01030201;
        8'h0A: out <= 32'h67A9CE67;
        8'h0B: out <= 32'h2B7D562B;
        8'h0C: out <= 32'hFE19E7FE;
        8'h0D: out <= 32'hD762B5D7;
        8'h0E: out <= 32'hABE64DAB;
        8'h0F: out <= 32'h769AEC76;
        8'h10: out <= 32'hCA458FCA;
        8'h11: out <= 32'h829D1F82;
        8'h12: out <= 32'hC94089C9;
        8'h13: out <= 32'h7D87FA7D;
        8'h14: out <= 32'hFA15EFFA;
        8'h15: out <= 32'h59EBB259;
        8'h16: out <= 32'h47C98E47;
        8'h17: out <= 32'hF00BFBF0;
        8'h18: out <= 32'hADEC41AD;
        8'h19: out <= 32'hD467B3D4;
        8'h1A: out <= 32'hA2FD5FA2;
        8'h1B: out <= 32'hAFEA45AF;
        8'h1C: out <= 32'h9CBF239C;
        8'h1D: out <= 32'hA4F753A4;
        8'h1E: out <= 32'h7296E472;
        8'h1F: out <= 32'hC05B9BC0;
        8'h20: out <= 32'hB7C275B7;
        8'h21: out <= 32'hFD1CE1FD;
        8'h22: out <= 32'h93AE3D93;
        8'h23: out <= 32'h266A4C26;
        8'h24: out <= 32'h365A6C36;
        8'h25: out <= 32'h3F417E3F;
        8'h26: out <= 32'hF702F5F7;
        8'h27: out <= 32'hCC4F83CC;
        8'h28: out <= 32'h345C6834;
        8'h29: out <= 32'hA5F451A5;
        8'h2A: out <= 32'hE534D1E5;
        8'h2B: out <= 32'hF108F9F1;
        8'h2C: out <= 32'h7193E271;
        8'h2D: out <= 32'hD873ABD8;
        8'h2E: out <= 32'h31536231;
        8'h2F: out <= 32'h153F2A15;
        8'h30: out <= 32'h040C0804;
        8'h31: out <= 32'hC75295C7;
        8'h32: out <= 32'h23654623;
        8'h33: out <= 32'hC35E9DC3;
        8'h34: out <= 32'h18283018;
        8'h35: out <= 32'h96A13796;
        8'h36: out <= 32'h050F0A05;
        8'h37: out <= 32'h9AB52F9A;
        8'h38: out <= 32'h07090E07;
        8'h39: out <= 32'h12362412;
        8'h3A: out <= 32'h809B1B80;
        8'h3B: out <= 32'hE23DDFE2;
        8'h3C: out <= 32'hEB26CDEB;
        8'h3D: out <= 32'h27694E27;
        8'h3E: out <= 32'hB2CD7FB2;
        8'h3F: out <= 32'h759FEA75;
        8'h40: out <= 32'h091B1209;
        8'h41: out <= 32'h839E1D83;
        8'h42: out <= 32'h2C74582C;
        8'h43: out <= 32'h1A2E341A;
        8'h44: out <= 32'h1B2D361B;
        8'h45: out <= 32'h6EB2DC6E;
        8'h46: out <= 32'h5AEEB45A;
        8'h47: out <= 32'hA0FB5BA0;
        8'h48: out <= 32'h52F6A452;
        8'h49: out <= 32'h3B4D763B;
        8'h4A: out <= 32'hD661B7D6;
        8'h4B: out <= 32'hB3CE7DB3;
        8'h4C: out <= 32'h297B5229;
        8'h4D: out <= 32'hE33EDDE3;
        8'h4E: out <= 32'h2F715E2F;
        8'h4F: out <= 32'h84971384;
        8'h50: out <= 32'h53F5A653;
        8'h51: out <= 32'hD168B9D1;
        8'h52: out <= 32'h00000000;
        8'h53: out <= 32'hED2CC1ED;
        8'h54: out <= 32'h20604020;
        8'h55: out <= 32'hFC1FE3FC;
        8'h56: out <= 32'hB1C879B1;
        8'h57: out <= 32'h5BEDB65B;
        8'h58: out <= 32'h6ABED46A;
        8'h59: out <= 32'hCB468DCB;
        8'h5A: out <= 32'hBED967BE;
        8'h5B: out <= 32'h394B7239;
        8'h5C: out <= 32'h4ADE944A;
        8'h5D: out <= 32'h4CD4984C;
        8'h5E: out <= 32'h58E8B058;
        8'h5F: out <= 32'hCF4A85CF;
        8'h60: out <= 32'hD06BBBD0;
        8'h61: out <= 32'hEF2AC5EF;
        8'h62: out <= 32'hAAE54FAA;
        8'h63: out <= 32'hFB16EDFB;
        8'h64: out <= 32'h43C58643;
        8'h65: out <= 32'h4DD79A4D;
        8'h66: out <= 32'h33556633;
        8'h67: out <= 32'h85941185;
        8'h68: out <= 32'h45CF8A45;
        8'h69: out <= 32'hF910E9F9;
        8'h6A: out <= 32'h02060402;
        8'h6B: out <= 32'h7F81FE7F;
        8'h6C: out <= 32'h50F0A050;
        8'h6D: out <= 32'h3C44783C;
        8'h6E: out <= 32'h9FBA259F;
        8'h6F: out <= 32'hA8E34BA8;
        8'h70: out <= 32'h51F3A251;
        8'h71: out <= 32'hA3FE5DA3;
        8'h72: out <= 32'h40C08040;
        8'h73: out <= 32'h8F8A058F;
        8'h74: out <= 32'h92AD3F92;
        8'h75: out <= 32'h9DBC219D;
        8'h76: out <= 32'h38487038;
        8'h77: out <= 32'hF504F1F5;
        8'h78: out <= 32'hBCDF63BC;
        8'h79: out <= 32'hB6C177B6;
        8'h7A: out <= 32'hDA75AFDA;
        8'h7B: out <= 32'h21634221;
        8'h7C: out <= 32'h10302010;
        8'h7D: out <= 32'hFF1AE5FF;
        8'h7E: out <= 32'hF30EFDF3;
        8'h7F: out <= 32'hD26DBFD2;
        8'h80: out <= 32'hCD4C81CD;
        8'h81: out <= 32'h0C14180C;
        8'h82: out <= 32'h13352613;
        8'h83: out <= 32'hEC2FC3EC;
        8'h84: out <= 32'h5FE1BE5F;
        8'h85: out <= 32'h97A23597;
        8'h86: out <= 32'h44CC8844;
        8'h87: out <= 32'h17392E17;
        8'h88: out <= 32'hC45793C4;
        8'h89: out <= 32'hA7F255A7;
        8'h8A: out <= 32'h7E82FC7E;
        8'h8B: out <= 32'h3D477A3D;
        8'h8C: out <= 32'h64ACC864;
        8'h8D: out <= 32'h5DE7BA5D;
        8'h8E: out <= 32'h192B3219;
        8'h8F: out <= 32'h7395E673;
        8'h90: out <= 32'h60A0C060;
        8'h91: out <= 32'h81981981;
        8'h92: out <= 32'h4FD19E4F;
        8'h93: out <= 32'hDC7FA3DC;
        8'h94: out <= 32'h22664422;
        8'h95: out <= 32'h2A7E542A;
        8'h96: out <= 32'h90AB3B90;
        8'h97: out <= 32'h88830B88;
        8'h98: out <= 32'h46CA8C46;
        8'h99: out <= 32'hEE29C7EE;
        8'h9A: out <= 32'hB8D36BB8;
        8'h9B: out <= 32'h143C2814;
        8'h9C: out <= 32'hDE79A7DE;
        8'h9D: out <= 32'h5EE2BC5E;
        8'h9E: out <= 32'h0B1D160B;
        8'h9F: out <= 32'hDB76ADDB;
        8'hA0: out <= 32'hE03BDBE0;
        8'hA1: out <= 32'h32566432;
        8'hA2: out <= 32'h3A4E743A;
        8'hA3: out <= 32'h0A1E140A;
        8'hA4: out <= 32'h49DB9249;
        8'hA5: out <= 32'h060A0C06;
        8'hA6: out <= 32'h246C4824;
        8'hA7: out <= 32'h5CE4B85C;
        8'hA8: out <= 32'hC25D9FC2;
        8'hA9: out <= 32'hD36EBDD3;
        8'hAA: out <= 32'hACEF43AC;
        8'hAB: out <= 32'h62A6C462;
        8'hAC: out <= 32'h91A83991;
        8'hAD: out <= 32'h95A43195;
        8'hAE: out <= 32'hE437D3E4;
        8'hAF: out <= 32'h798BF279;
        8'hB0: out <= 32'hE732D5E7;
        8'hB1: out <= 32'hC8438BC8;
        8'hB2: out <= 32'h37596E37;
        8'hB3: out <= 32'h6DB7DA6D;
        8'hB4: out <= 32'h8D8C018D;
        8'hB5: out <= 32'hD564B1D5;
        8'hB6: out <= 32'h4ED29C4E;
        8'hB7: out <= 32'hA9E049A9;
        8'hB8: out <= 32'h6CB4D86C;
        8'hB9: out <= 32'h56FAAC56;
        8'hBA: out <= 32'hF407F3F4;
        8'hBB: out <= 32'hEA25CFEA;
        8'hBC: out <= 32'h65AFCA65;
        8'hBD: out <= 32'h7A8EF47A;
        8'hBE: out <= 32'hAEE947AE;
        8'hBF: out <= 32'h08181008;
        8'hC0: out <= 32'hBAD56FBA;
        8'hC1: out <= 32'h7888F078;
        8'hC2: out <= 32'h256F4A25;
        8'hC3: out <= 32'h2E725C2E;
        8'hC4: out <= 32'h1C24381C;
        8'hC5: out <= 32'hA6F157A6;
        8'hC6: out <= 32'hB4C773B4;
        8'hC7: out <= 32'hC65197C6;
        8'hC8: out <= 32'hE823CBE8;
        8'hC9: out <= 32'hDD7CA1DD;
        8'hCA: out <= 32'h749CE874;
        8'hCB: out <= 32'h1F213E1F;
        8'hCC: out <= 32'h4BDD964B;
        8'hCD: out <= 32'hBDDC61BD;
        8'hCE: out <= 32'h8B860D8B;
        8'hCF: out <= 32'h8A850F8A;
        8'hD0: out <= 32'h7090E070;
        8'hD1: out <= 32'h3E427C3E;
        8'hD2: out <= 32'hB5C471B5;
        8'hD3: out <= 32'h66AACC66;
        8'hD4: out <= 32'h48D89048;
        8'hD5: out <= 32'h03050603;
        8'hD6: out <= 32'hF601F7F6;
        8'hD7: out <= 32'h0E121C0E;
        8'hD8: out <= 32'h61A3C261;
        8'hD9: out <= 32'h355F6A35;
        8'hDA: out <= 32'h57F9AE57;
        8'hDB: out <= 32'hB9D069B9;
        8'hDC: out <= 32'h86911786;
        8'hDD: out <= 32'hC15899C1;
        8'hDE: out <= 32'h1D273A1D;
        8'hDF: out <= 32'h9EB9279E;
        8'hE0: out <= 32'hE138D9E1;
        8'hE1: out <= 32'hF813EBF8;
        8'hE2: out <= 32'h98B32B98;
        8'hE3: out <= 32'h11332211;
        8'hE4: out <= 32'h69BBD269;
        8'hE5: out <= 32'hD970A9D9;
        8'hE6: out <= 32'h8E89078E;
        8'hE7: out <= 32'h94A73394;
        8'hE8: out <= 32'h9BB62D9B;
        8'hE9: out <= 32'h1E223C1E;
        8'hEA: out <= 32'h87921587;
        8'hEB: out <= 32'hE920C9E9;
        8'hEC: out <= 32'hCE4987CE;
        8'hED: out <= 32'h55FFAA55;
        8'hEE: out <= 32'h28785028;
        8'hEF: out <= 32'hDF7AA5DF;
        8'hF0: out <= 32'h8C8F038C;
        8'hF1: out <= 32'hA1F859A1;
        8'hF2: out <= 32'h89800989;
        8'hF3: out <= 32'h0D171A0D;
        8'hF4: out <= 32'hBFDA65BF;
        8'hF5: out <= 32'hE631D7E6;
        8'hF6: out <= 32'h42C68442;
        8'hF7: out <= 32'h68B8D068;
        8'hF8: out <= 32'h41C38241;
        8'hF9: out <= 32'h99B02999;
        8'hFA: out <= 32'h2D775A2D;
        8'hFB: out <= 32'h0F111E0F;
        8'hFC: out <= 32'hB0CB7BB0;
        8'hFD: out <= 32'h54FCA854;
        8'hFE: out <= 32'hBBD66DBB;
        8'hFF: out <= 32'h163A2C16;
        endcase
    end
endmodule
