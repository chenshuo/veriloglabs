../basic/Rcon.sv