../sbox/key_schedule.sv