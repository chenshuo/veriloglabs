module Te0box(in, clk, out);
    input [7:0] in;
    input clk;
    output[31:0] out;

    reg[31:0] out;

    always @(posedge clk)
    begin
        case (in)
        8'h00: out <= 32'hC66363A5;
        8'h01: out <= 32'hF87C7C84;
        8'h02: out <= 32'hEE777799;
        8'h03: out <= 32'hF67B7B8D;
        8'h04: out <= 32'hFFF2F20D;
        8'h05: out <= 32'hD66B6BBD;
        8'h06: out <= 32'hDE6F6FB1;
        8'h07: out <= 32'h91C5C554;
        8'h08: out <= 32'h60303050;
        8'h09: out <= 32'h02010103;
        8'h0A: out <= 32'hCE6767A9;
        8'h0B: out <= 32'h562B2B7D;
        8'h0C: out <= 32'hE7FEFE19;
        8'h0D: out <= 32'hB5D7D762;
        8'h0E: out <= 32'h4DABABE6;
        8'h0F: out <= 32'hEC76769A;
        8'h10: out <= 32'h8FCACA45;
        8'h11: out <= 32'h1F82829D;
        8'h12: out <= 32'h89C9C940;
        8'h13: out <= 32'hFA7D7D87;
        8'h14: out <= 32'hEFFAFA15;
        8'h15: out <= 32'hB25959EB;
        8'h16: out <= 32'h8E4747C9;
        8'h17: out <= 32'hFBF0F00B;
        8'h18: out <= 32'h41ADADEC;
        8'h19: out <= 32'hB3D4D467;
        8'h1A: out <= 32'h5FA2A2FD;
        8'h1B: out <= 32'h45AFAFEA;
        8'h1C: out <= 32'h239C9CBF;
        8'h1D: out <= 32'h53A4A4F7;
        8'h1E: out <= 32'hE4727296;
        8'h1F: out <= 32'h9BC0C05B;
        8'h20: out <= 32'h75B7B7C2;
        8'h21: out <= 32'hE1FDFD1C;
        8'h22: out <= 32'h3D9393AE;
        8'h23: out <= 32'h4C26266A;
        8'h24: out <= 32'h6C36365A;
        8'h25: out <= 32'h7E3F3F41;
        8'h26: out <= 32'hF5F7F702;
        8'h27: out <= 32'h83CCCC4F;
        8'h28: out <= 32'h6834345C;
        8'h29: out <= 32'h51A5A5F4;
        8'h2A: out <= 32'hD1E5E534;
        8'h2B: out <= 32'hF9F1F108;
        8'h2C: out <= 32'hE2717193;
        8'h2D: out <= 32'hABD8D873;
        8'h2E: out <= 32'h62313153;
        8'h2F: out <= 32'h2A15153F;
        8'h30: out <= 32'h0804040C;
        8'h31: out <= 32'h95C7C752;
        8'h32: out <= 32'h46232365;
        8'h33: out <= 32'h9DC3C35E;
        8'h34: out <= 32'h30181828;
        8'h35: out <= 32'h379696A1;
        8'h36: out <= 32'h0A05050F;
        8'h37: out <= 32'h2F9A9AB5;
        8'h38: out <= 32'h0E070709;
        8'h39: out <= 32'h24121236;
        8'h3A: out <= 32'h1B80809B;
        8'h3B: out <= 32'hDFE2E23D;
        8'h3C: out <= 32'hCDEBEB26;
        8'h3D: out <= 32'h4E272769;
        8'h3E: out <= 32'h7FB2B2CD;
        8'h3F: out <= 32'hEA75759F;
        8'h40: out <= 32'h1209091B;
        8'h41: out <= 32'h1D83839E;
        8'h42: out <= 32'h582C2C74;
        8'h43: out <= 32'h341A1A2E;
        8'h44: out <= 32'h361B1B2D;
        8'h45: out <= 32'hDC6E6EB2;
        8'h46: out <= 32'hB45A5AEE;
        8'h47: out <= 32'h5BA0A0FB;
        8'h48: out <= 32'hA45252F6;
        8'h49: out <= 32'h763B3B4D;
        8'h4A: out <= 32'hB7D6D661;
        8'h4B: out <= 32'h7DB3B3CE;
        8'h4C: out <= 32'h5229297B;
        8'h4D: out <= 32'hDDE3E33E;
        8'h4E: out <= 32'h5E2F2F71;
        8'h4F: out <= 32'h13848497;
        8'h50: out <= 32'hA65353F5;
        8'h51: out <= 32'hB9D1D168;
        8'h52: out <= 32'h00000000;
        8'h53: out <= 32'hC1EDED2C;
        8'h54: out <= 32'h40202060;
        8'h55: out <= 32'hE3FCFC1F;
        8'h56: out <= 32'h79B1B1C8;
        8'h57: out <= 32'hB65B5BED;
        8'h58: out <= 32'hD46A6ABE;
        8'h59: out <= 32'h8DCBCB46;
        8'h5A: out <= 32'h67BEBED9;
        8'h5B: out <= 32'h7239394B;
        8'h5C: out <= 32'h944A4ADE;
        8'h5D: out <= 32'h984C4CD4;
        8'h5E: out <= 32'hB05858E8;
        8'h5F: out <= 32'h85CFCF4A;
        8'h60: out <= 32'hBBD0D06B;
        8'h61: out <= 32'hC5EFEF2A;
        8'h62: out <= 32'h4FAAAAE5;
        8'h63: out <= 32'hEDFBFB16;
        8'h64: out <= 32'h864343C5;
        8'h65: out <= 32'h9A4D4DD7;
        8'h66: out <= 32'h66333355;
        8'h67: out <= 32'h11858594;
        8'h68: out <= 32'h8A4545CF;
        8'h69: out <= 32'hE9F9F910;
        8'h6A: out <= 32'h04020206;
        8'h6B: out <= 32'hFE7F7F81;
        8'h6C: out <= 32'hA05050F0;
        8'h6D: out <= 32'h783C3C44;
        8'h6E: out <= 32'h259F9FBA;
        8'h6F: out <= 32'h4BA8A8E3;
        8'h70: out <= 32'hA25151F3;
        8'h71: out <= 32'h5DA3A3FE;
        8'h72: out <= 32'h804040C0;
        8'h73: out <= 32'h058F8F8A;
        8'h74: out <= 32'h3F9292AD;
        8'h75: out <= 32'h219D9DBC;
        8'h76: out <= 32'h70383848;
        8'h77: out <= 32'hF1F5F504;
        8'h78: out <= 32'h63BCBCDF;
        8'h79: out <= 32'h77B6B6C1;
        8'h7A: out <= 32'hAFDADA75;
        8'h7B: out <= 32'h42212163;
        8'h7C: out <= 32'h20101030;
        8'h7D: out <= 32'hE5FFFF1A;
        8'h7E: out <= 32'hFDF3F30E;
        8'h7F: out <= 32'hBFD2D26D;
        8'h80: out <= 32'h81CDCD4C;
        8'h81: out <= 32'h180C0C14;
        8'h82: out <= 32'h26131335;
        8'h83: out <= 32'hC3ECEC2F;
        8'h84: out <= 32'hBE5F5FE1;
        8'h85: out <= 32'h359797A2;
        8'h86: out <= 32'h884444CC;
        8'h87: out <= 32'h2E171739;
        8'h88: out <= 32'h93C4C457;
        8'h89: out <= 32'h55A7A7F2;
        8'h8A: out <= 32'hFC7E7E82;
        8'h8B: out <= 32'h7A3D3D47;
        8'h8C: out <= 32'hC86464AC;
        8'h8D: out <= 32'hBA5D5DE7;
        8'h8E: out <= 32'h3219192B;
        8'h8F: out <= 32'hE6737395;
        8'h90: out <= 32'hC06060A0;
        8'h91: out <= 32'h19818198;
        8'h92: out <= 32'h9E4F4FD1;
        8'h93: out <= 32'hA3DCDC7F;
        8'h94: out <= 32'h44222266;
        8'h95: out <= 32'h542A2A7E;
        8'h96: out <= 32'h3B9090AB;
        8'h97: out <= 32'h0B888883;
        8'h98: out <= 32'h8C4646CA;
        8'h99: out <= 32'hC7EEEE29;
        8'h9A: out <= 32'h6BB8B8D3;
        8'h9B: out <= 32'h2814143C;
        8'h9C: out <= 32'hA7DEDE79;
        8'h9D: out <= 32'hBC5E5EE2;
        8'h9E: out <= 32'h160B0B1D;
        8'h9F: out <= 32'hADDBDB76;
        8'hA0: out <= 32'hDBE0E03B;
        8'hA1: out <= 32'h64323256;
        8'hA2: out <= 32'h743A3A4E;
        8'hA3: out <= 32'h140A0A1E;
        8'hA4: out <= 32'h924949DB;
        8'hA5: out <= 32'h0C06060A;
        8'hA6: out <= 32'h4824246C;
        8'hA7: out <= 32'hB85C5CE4;
        8'hA8: out <= 32'h9FC2C25D;
        8'hA9: out <= 32'hBDD3D36E;
        8'hAA: out <= 32'h43ACACEF;
        8'hAB: out <= 32'hC46262A6;
        8'hAC: out <= 32'h399191A8;
        8'hAD: out <= 32'h319595A4;
        8'hAE: out <= 32'hD3E4E437;
        8'hAF: out <= 32'hF279798B;
        8'hB0: out <= 32'hD5E7E732;
        8'hB1: out <= 32'h8BC8C843;
        8'hB2: out <= 32'h6E373759;
        8'hB3: out <= 32'hDA6D6DB7;
        8'hB4: out <= 32'h018D8D8C;
        8'hB5: out <= 32'hB1D5D564;
        8'hB6: out <= 32'h9C4E4ED2;
        8'hB7: out <= 32'h49A9A9E0;
        8'hB8: out <= 32'hD86C6CB4;
        8'hB9: out <= 32'hAC5656FA;
        8'hBA: out <= 32'hF3F4F407;
        8'hBB: out <= 32'hCFEAEA25;
        8'hBC: out <= 32'hCA6565AF;
        8'hBD: out <= 32'hF47A7A8E;
        8'hBE: out <= 32'h47AEAEE9;
        8'hBF: out <= 32'h10080818;
        8'hC0: out <= 32'h6FBABAD5;
        8'hC1: out <= 32'hF0787888;
        8'hC2: out <= 32'h4A25256F;
        8'hC3: out <= 32'h5C2E2E72;
        8'hC4: out <= 32'h381C1C24;
        8'hC5: out <= 32'h57A6A6F1;
        8'hC6: out <= 32'h73B4B4C7;
        8'hC7: out <= 32'h97C6C651;
        8'hC8: out <= 32'hCBE8E823;
        8'hC9: out <= 32'hA1DDDD7C;
        8'hCA: out <= 32'hE874749C;
        8'hCB: out <= 32'h3E1F1F21;
        8'hCC: out <= 32'h964B4BDD;
        8'hCD: out <= 32'h61BDBDDC;
        8'hCE: out <= 32'h0D8B8B86;
        8'hCF: out <= 32'h0F8A8A85;
        8'hD0: out <= 32'hE0707090;
        8'hD1: out <= 32'h7C3E3E42;
        8'hD2: out <= 32'h71B5B5C4;
        8'hD3: out <= 32'hCC6666AA;
        8'hD4: out <= 32'h904848D8;
        8'hD5: out <= 32'h06030305;
        8'hD6: out <= 32'hF7F6F601;
        8'hD7: out <= 32'h1C0E0E12;
        8'hD8: out <= 32'hC26161A3;
        8'hD9: out <= 32'h6A35355F;
        8'hDA: out <= 32'hAE5757F9;
        8'hDB: out <= 32'h69B9B9D0;
        8'hDC: out <= 32'h17868691;
        8'hDD: out <= 32'h99C1C158;
        8'hDE: out <= 32'h3A1D1D27;
        8'hDF: out <= 32'h279E9EB9;
        8'hE0: out <= 32'hD9E1E138;
        8'hE1: out <= 32'hEBF8F813;
        8'hE2: out <= 32'h2B9898B3;
        8'hE3: out <= 32'h22111133;
        8'hE4: out <= 32'hD26969BB;
        8'hE5: out <= 32'hA9D9D970;
        8'hE6: out <= 32'h078E8E89;
        8'hE7: out <= 32'h339494A7;
        8'hE8: out <= 32'h2D9B9BB6;
        8'hE9: out <= 32'h3C1E1E22;
        8'hEA: out <= 32'h15878792;
        8'hEB: out <= 32'hC9E9E920;
        8'hEC: out <= 32'h87CECE49;
        8'hED: out <= 32'hAA5555FF;
        8'hEE: out <= 32'h50282878;
        8'hEF: out <= 32'hA5DFDF7A;
        8'hF0: out <= 32'h038C8C8F;
        8'hF1: out <= 32'h59A1A1F8;
        8'hF2: out <= 32'h09898980;
        8'hF3: out <= 32'h1A0D0D17;
        8'hF4: out <= 32'h65BFBFDA;
        8'hF5: out <= 32'hD7E6E631;
        8'hF6: out <= 32'h844242C6;
        8'hF7: out <= 32'hD06868B8;
        8'hF8: out <= 32'h824141C3;
        8'hF9: out <= 32'h299999B0;
        8'hFA: out <= 32'h5A2D2D77;
        8'hFB: out <= 32'h1E0F0F11;
        8'hFC: out <= 32'h7BB0B0CB;
        8'hFD: out <= 32'hA85454FC;
        8'hFE: out <= 32'h6DBBBBD6;
        8'hFF: out <= 32'h2C16163A;
        endcase
    end
endmodule
