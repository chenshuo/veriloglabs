module Te1box(in, clk, out);
    input [7:0] in;
    input clk;
    output[31:0] out;

    reg[31:0] out;

    always @(posedge clk)
    begin
        case (in)
        8'h00: out <= 32'hA5C66363;
        8'h01: out <= 32'h84F87C7C;
        8'h02: out <= 32'h99EE7777;
        8'h03: out <= 32'h8DF67B7B;
        8'h04: out <= 32'h0DFFF2F2;
        8'h05: out <= 32'hBDD66B6B;
        8'h06: out <= 32'hB1DE6F6F;
        8'h07: out <= 32'h5491C5C5;
        8'h08: out <= 32'h50603030;
        8'h09: out <= 32'h03020101;
        8'h0A: out <= 32'hA9CE6767;
        8'h0B: out <= 32'h7D562B2B;
        8'h0C: out <= 32'h19E7FEFE;
        8'h0D: out <= 32'h62B5D7D7;
        8'h0E: out <= 32'hE64DABAB;
        8'h0F: out <= 32'h9AEC7676;
        8'h10: out <= 32'h458FCACA;
        8'h11: out <= 32'h9D1F8282;
        8'h12: out <= 32'h4089C9C9;
        8'h13: out <= 32'h87FA7D7D;
        8'h14: out <= 32'h15EFFAFA;
        8'h15: out <= 32'hEBB25959;
        8'h16: out <= 32'hC98E4747;
        8'h17: out <= 32'h0BFBF0F0;
        8'h18: out <= 32'hEC41ADAD;
        8'h19: out <= 32'h67B3D4D4;
        8'h1A: out <= 32'hFD5FA2A2;
        8'h1B: out <= 32'hEA45AFAF;
        8'h1C: out <= 32'hBF239C9C;
        8'h1D: out <= 32'hF753A4A4;
        8'h1E: out <= 32'h96E47272;
        8'h1F: out <= 32'h5B9BC0C0;
        8'h20: out <= 32'hC275B7B7;
        8'h21: out <= 32'h1CE1FDFD;
        8'h22: out <= 32'hAE3D9393;
        8'h23: out <= 32'h6A4C2626;
        8'h24: out <= 32'h5A6C3636;
        8'h25: out <= 32'h417E3F3F;
        8'h26: out <= 32'h02F5F7F7;
        8'h27: out <= 32'h4F83CCCC;
        8'h28: out <= 32'h5C683434;
        8'h29: out <= 32'hF451A5A5;
        8'h2A: out <= 32'h34D1E5E5;
        8'h2B: out <= 32'h08F9F1F1;
        8'h2C: out <= 32'h93E27171;
        8'h2D: out <= 32'h73ABD8D8;
        8'h2E: out <= 32'h53623131;
        8'h2F: out <= 32'h3F2A1515;
        8'h30: out <= 32'h0C080404;
        8'h31: out <= 32'h5295C7C7;
        8'h32: out <= 32'h65462323;
        8'h33: out <= 32'h5E9DC3C3;
        8'h34: out <= 32'h28301818;
        8'h35: out <= 32'hA1379696;
        8'h36: out <= 32'h0F0A0505;
        8'h37: out <= 32'hB52F9A9A;
        8'h38: out <= 32'h090E0707;
        8'h39: out <= 32'h36241212;
        8'h3A: out <= 32'h9B1B8080;
        8'h3B: out <= 32'h3DDFE2E2;
        8'h3C: out <= 32'h26CDEBEB;
        8'h3D: out <= 32'h694E2727;
        8'h3E: out <= 32'hCD7FB2B2;
        8'h3F: out <= 32'h9FEA7575;
        8'h40: out <= 32'h1B120909;
        8'h41: out <= 32'h9E1D8383;
        8'h42: out <= 32'h74582C2C;
        8'h43: out <= 32'h2E341A1A;
        8'h44: out <= 32'h2D361B1B;
        8'h45: out <= 32'hB2DC6E6E;
        8'h46: out <= 32'hEEB45A5A;
        8'h47: out <= 32'hFB5BA0A0;
        8'h48: out <= 32'hF6A45252;
        8'h49: out <= 32'h4D763B3B;
        8'h4A: out <= 32'h61B7D6D6;
        8'h4B: out <= 32'hCE7DB3B3;
        8'h4C: out <= 32'h7B522929;
        8'h4D: out <= 32'h3EDDE3E3;
        8'h4E: out <= 32'h715E2F2F;
        8'h4F: out <= 32'h97138484;
        8'h50: out <= 32'hF5A65353;
        8'h51: out <= 32'h68B9D1D1;
        8'h52: out <= 32'h00000000;
        8'h53: out <= 32'h2CC1EDED;
        8'h54: out <= 32'h60402020;
        8'h55: out <= 32'h1FE3FCFC;
        8'h56: out <= 32'hC879B1B1;
        8'h57: out <= 32'hEDB65B5B;
        8'h58: out <= 32'hBED46A6A;
        8'h59: out <= 32'h468DCBCB;
        8'h5A: out <= 32'hD967BEBE;
        8'h5B: out <= 32'h4B723939;
        8'h5C: out <= 32'hDE944A4A;
        8'h5D: out <= 32'hD4984C4C;
        8'h5E: out <= 32'hE8B05858;
        8'h5F: out <= 32'h4A85CFCF;
        8'h60: out <= 32'h6BBBD0D0;
        8'h61: out <= 32'h2AC5EFEF;
        8'h62: out <= 32'hE54FAAAA;
        8'h63: out <= 32'h16EDFBFB;
        8'h64: out <= 32'hC5864343;
        8'h65: out <= 32'hD79A4D4D;
        8'h66: out <= 32'h55663333;
        8'h67: out <= 32'h94118585;
        8'h68: out <= 32'hCF8A4545;
        8'h69: out <= 32'h10E9F9F9;
        8'h6A: out <= 32'h06040202;
        8'h6B: out <= 32'h81FE7F7F;
        8'h6C: out <= 32'hF0A05050;
        8'h6D: out <= 32'h44783C3C;
        8'h6E: out <= 32'hBA259F9F;
        8'h6F: out <= 32'hE34BA8A8;
        8'h70: out <= 32'hF3A25151;
        8'h71: out <= 32'hFE5DA3A3;
        8'h72: out <= 32'hC0804040;
        8'h73: out <= 32'h8A058F8F;
        8'h74: out <= 32'hAD3F9292;
        8'h75: out <= 32'hBC219D9D;
        8'h76: out <= 32'h48703838;
        8'h77: out <= 32'h04F1F5F5;
        8'h78: out <= 32'hDF63BCBC;
        8'h79: out <= 32'hC177B6B6;
        8'h7A: out <= 32'h75AFDADA;
        8'h7B: out <= 32'h63422121;
        8'h7C: out <= 32'h30201010;
        8'h7D: out <= 32'h1AE5FFFF;
        8'h7E: out <= 32'h0EFDF3F3;
        8'h7F: out <= 32'h6DBFD2D2;
        8'h80: out <= 32'h4C81CDCD;
        8'h81: out <= 32'h14180C0C;
        8'h82: out <= 32'h35261313;
        8'h83: out <= 32'h2FC3ECEC;
        8'h84: out <= 32'hE1BE5F5F;
        8'h85: out <= 32'hA2359797;
        8'h86: out <= 32'hCC884444;
        8'h87: out <= 32'h392E1717;
        8'h88: out <= 32'h5793C4C4;
        8'h89: out <= 32'hF255A7A7;
        8'h8A: out <= 32'h82FC7E7E;
        8'h8B: out <= 32'h477A3D3D;
        8'h8C: out <= 32'hACC86464;
        8'h8D: out <= 32'hE7BA5D5D;
        8'h8E: out <= 32'h2B321919;
        8'h8F: out <= 32'h95E67373;
        8'h90: out <= 32'hA0C06060;
        8'h91: out <= 32'h98198181;
        8'h92: out <= 32'hD19E4F4F;
        8'h93: out <= 32'h7FA3DCDC;
        8'h94: out <= 32'h66442222;
        8'h95: out <= 32'h7E542A2A;
        8'h96: out <= 32'hAB3B9090;
        8'h97: out <= 32'h830B8888;
        8'h98: out <= 32'hCA8C4646;
        8'h99: out <= 32'h29C7EEEE;
        8'h9A: out <= 32'hD36BB8B8;
        8'h9B: out <= 32'h3C281414;
        8'h9C: out <= 32'h79A7DEDE;
        8'h9D: out <= 32'hE2BC5E5E;
        8'h9E: out <= 32'h1D160B0B;
        8'h9F: out <= 32'h76ADDBDB;
        8'hA0: out <= 32'h3BDBE0E0;
        8'hA1: out <= 32'h56643232;
        8'hA2: out <= 32'h4E743A3A;
        8'hA3: out <= 32'h1E140A0A;
        8'hA4: out <= 32'hDB924949;
        8'hA5: out <= 32'h0A0C0606;
        8'hA6: out <= 32'h6C482424;
        8'hA7: out <= 32'hE4B85C5C;
        8'hA8: out <= 32'h5D9FC2C2;
        8'hA9: out <= 32'h6EBDD3D3;
        8'hAA: out <= 32'hEF43ACAC;
        8'hAB: out <= 32'hA6C46262;
        8'hAC: out <= 32'hA8399191;
        8'hAD: out <= 32'hA4319595;
        8'hAE: out <= 32'h37D3E4E4;
        8'hAF: out <= 32'h8BF27979;
        8'hB0: out <= 32'h32D5E7E7;
        8'hB1: out <= 32'h438BC8C8;
        8'hB2: out <= 32'h596E3737;
        8'hB3: out <= 32'hB7DA6D6D;
        8'hB4: out <= 32'h8C018D8D;
        8'hB5: out <= 32'h64B1D5D5;
        8'hB6: out <= 32'hD29C4E4E;
        8'hB7: out <= 32'hE049A9A9;
        8'hB8: out <= 32'hB4D86C6C;
        8'hB9: out <= 32'hFAAC5656;
        8'hBA: out <= 32'h07F3F4F4;
        8'hBB: out <= 32'h25CFEAEA;
        8'hBC: out <= 32'hAFCA6565;
        8'hBD: out <= 32'h8EF47A7A;
        8'hBE: out <= 32'hE947AEAE;
        8'hBF: out <= 32'h18100808;
        8'hC0: out <= 32'hD56FBABA;
        8'hC1: out <= 32'h88F07878;
        8'hC2: out <= 32'h6F4A2525;
        8'hC3: out <= 32'h725C2E2E;
        8'hC4: out <= 32'h24381C1C;
        8'hC5: out <= 32'hF157A6A6;
        8'hC6: out <= 32'hC773B4B4;
        8'hC7: out <= 32'h5197C6C6;
        8'hC8: out <= 32'h23CBE8E8;
        8'hC9: out <= 32'h7CA1DDDD;
        8'hCA: out <= 32'h9CE87474;
        8'hCB: out <= 32'h213E1F1F;
        8'hCC: out <= 32'hDD964B4B;
        8'hCD: out <= 32'hDC61BDBD;
        8'hCE: out <= 32'h860D8B8B;
        8'hCF: out <= 32'h850F8A8A;
        8'hD0: out <= 32'h90E07070;
        8'hD1: out <= 32'h427C3E3E;
        8'hD2: out <= 32'hC471B5B5;
        8'hD3: out <= 32'hAACC6666;
        8'hD4: out <= 32'hD8904848;
        8'hD5: out <= 32'h05060303;
        8'hD6: out <= 32'h01F7F6F6;
        8'hD7: out <= 32'h121C0E0E;
        8'hD8: out <= 32'hA3C26161;
        8'hD9: out <= 32'h5F6A3535;
        8'hDA: out <= 32'hF9AE5757;
        8'hDB: out <= 32'hD069B9B9;
        8'hDC: out <= 32'h91178686;
        8'hDD: out <= 32'h5899C1C1;
        8'hDE: out <= 32'h273A1D1D;
        8'hDF: out <= 32'hB9279E9E;
        8'hE0: out <= 32'h38D9E1E1;
        8'hE1: out <= 32'h13EBF8F8;
        8'hE2: out <= 32'hB32B9898;
        8'hE3: out <= 32'h33221111;
        8'hE4: out <= 32'hBBD26969;
        8'hE5: out <= 32'h70A9D9D9;
        8'hE6: out <= 32'h89078E8E;
        8'hE7: out <= 32'hA7339494;
        8'hE8: out <= 32'hB62D9B9B;
        8'hE9: out <= 32'h223C1E1E;
        8'hEA: out <= 32'h92158787;
        8'hEB: out <= 32'h20C9E9E9;
        8'hEC: out <= 32'h4987CECE;
        8'hED: out <= 32'hFFAA5555;
        8'hEE: out <= 32'h78502828;
        8'hEF: out <= 32'h7AA5DFDF;
        8'hF0: out <= 32'h8F038C8C;
        8'hF1: out <= 32'hF859A1A1;
        8'hF2: out <= 32'h80098989;
        8'hF3: out <= 32'h171A0D0D;
        8'hF4: out <= 32'hDA65BFBF;
        8'hF5: out <= 32'h31D7E6E6;
        8'hF6: out <= 32'hC6844242;
        8'hF7: out <= 32'hB8D06868;
        8'hF8: out <= 32'hC3824141;
        8'hF9: out <= 32'hB0299999;
        8'hFA: out <= 32'h775A2D2D;
        8'hFB: out <= 32'h111E0F0F;
        8'hFC: out <= 32'hCB7BB0B0;
        8'hFD: out <= 32'hFCA85454;
        8'hFE: out <= 32'hD66DBBBB;
        8'hFF: out <= 32'h3A2C1616;
        endcase
    end
endmodule
