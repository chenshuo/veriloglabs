../sbox/Rcon.sv