../sbox/Sbox.sv