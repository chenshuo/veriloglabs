../tbox/aes_encrypt_core_tb.sv