../tboxdp/Tbox.sv