module Te3box(in, clk, out);
    input [7:0] in;
    input clk;
    output[31:0] out;

    reg[31:0] out;

    always @(posedge clk)
    begin
        case (in)
        8'h00: out <= 32'h6363A5C6;
        8'h01: out <= 32'h7C7C84F8;
        8'h02: out <= 32'h777799EE;
        8'h03: out <= 32'h7B7B8DF6;
        8'h04: out <= 32'hF2F20DFF;
        8'h05: out <= 32'h6B6BBDD6;
        8'h06: out <= 32'h6F6FB1DE;
        8'h07: out <= 32'hC5C55491;
        8'h08: out <= 32'h30305060;
        8'h09: out <= 32'h01010302;
        8'h0A: out <= 32'h6767A9CE;
        8'h0B: out <= 32'h2B2B7D56;
        8'h0C: out <= 32'hFEFE19E7;
        8'h0D: out <= 32'hD7D762B5;
        8'h0E: out <= 32'hABABE64D;
        8'h0F: out <= 32'h76769AEC;
        8'h10: out <= 32'hCACA458F;
        8'h11: out <= 32'h82829D1F;
        8'h12: out <= 32'hC9C94089;
        8'h13: out <= 32'h7D7D87FA;
        8'h14: out <= 32'hFAFA15EF;
        8'h15: out <= 32'h5959EBB2;
        8'h16: out <= 32'h4747C98E;
        8'h17: out <= 32'hF0F00BFB;
        8'h18: out <= 32'hADADEC41;
        8'h19: out <= 32'hD4D467B3;
        8'h1A: out <= 32'hA2A2FD5F;
        8'h1B: out <= 32'hAFAFEA45;
        8'h1C: out <= 32'h9C9CBF23;
        8'h1D: out <= 32'hA4A4F753;
        8'h1E: out <= 32'h727296E4;
        8'h1F: out <= 32'hC0C05B9B;
        8'h20: out <= 32'hB7B7C275;
        8'h21: out <= 32'hFDFD1CE1;
        8'h22: out <= 32'h9393AE3D;
        8'h23: out <= 32'h26266A4C;
        8'h24: out <= 32'h36365A6C;
        8'h25: out <= 32'h3F3F417E;
        8'h26: out <= 32'hF7F702F5;
        8'h27: out <= 32'hCCCC4F83;
        8'h28: out <= 32'h34345C68;
        8'h29: out <= 32'hA5A5F451;
        8'h2A: out <= 32'hE5E534D1;
        8'h2B: out <= 32'hF1F108F9;
        8'h2C: out <= 32'h717193E2;
        8'h2D: out <= 32'hD8D873AB;
        8'h2E: out <= 32'h31315362;
        8'h2F: out <= 32'h15153F2A;
        8'h30: out <= 32'h04040C08;
        8'h31: out <= 32'hC7C75295;
        8'h32: out <= 32'h23236546;
        8'h33: out <= 32'hC3C35E9D;
        8'h34: out <= 32'h18182830;
        8'h35: out <= 32'h9696A137;
        8'h36: out <= 32'h05050F0A;
        8'h37: out <= 32'h9A9AB52F;
        8'h38: out <= 32'h0707090E;
        8'h39: out <= 32'h12123624;
        8'h3A: out <= 32'h80809B1B;
        8'h3B: out <= 32'hE2E23DDF;
        8'h3C: out <= 32'hEBEB26CD;
        8'h3D: out <= 32'h2727694E;
        8'h3E: out <= 32'hB2B2CD7F;
        8'h3F: out <= 32'h75759FEA;
        8'h40: out <= 32'h09091B12;
        8'h41: out <= 32'h83839E1D;
        8'h42: out <= 32'h2C2C7458;
        8'h43: out <= 32'h1A1A2E34;
        8'h44: out <= 32'h1B1B2D36;
        8'h45: out <= 32'h6E6EB2DC;
        8'h46: out <= 32'h5A5AEEB4;
        8'h47: out <= 32'hA0A0FB5B;
        8'h48: out <= 32'h5252F6A4;
        8'h49: out <= 32'h3B3B4D76;
        8'h4A: out <= 32'hD6D661B7;
        8'h4B: out <= 32'hB3B3CE7D;
        8'h4C: out <= 32'h29297B52;
        8'h4D: out <= 32'hE3E33EDD;
        8'h4E: out <= 32'h2F2F715E;
        8'h4F: out <= 32'h84849713;
        8'h50: out <= 32'h5353F5A6;
        8'h51: out <= 32'hD1D168B9;
        8'h52: out <= 32'h00000000;
        8'h53: out <= 32'hEDED2CC1;
        8'h54: out <= 32'h20206040;
        8'h55: out <= 32'hFCFC1FE3;
        8'h56: out <= 32'hB1B1C879;
        8'h57: out <= 32'h5B5BEDB6;
        8'h58: out <= 32'h6A6ABED4;
        8'h59: out <= 32'hCBCB468D;
        8'h5A: out <= 32'hBEBED967;
        8'h5B: out <= 32'h39394B72;
        8'h5C: out <= 32'h4A4ADE94;
        8'h5D: out <= 32'h4C4CD498;
        8'h5E: out <= 32'h5858E8B0;
        8'h5F: out <= 32'hCFCF4A85;
        8'h60: out <= 32'hD0D06BBB;
        8'h61: out <= 32'hEFEF2AC5;
        8'h62: out <= 32'hAAAAE54F;
        8'h63: out <= 32'hFBFB16ED;
        8'h64: out <= 32'h4343C586;
        8'h65: out <= 32'h4D4DD79A;
        8'h66: out <= 32'h33335566;
        8'h67: out <= 32'h85859411;
        8'h68: out <= 32'h4545CF8A;
        8'h69: out <= 32'hF9F910E9;
        8'h6A: out <= 32'h02020604;
        8'h6B: out <= 32'h7F7F81FE;
        8'h6C: out <= 32'h5050F0A0;
        8'h6D: out <= 32'h3C3C4478;
        8'h6E: out <= 32'h9F9FBA25;
        8'h6F: out <= 32'hA8A8E34B;
        8'h70: out <= 32'h5151F3A2;
        8'h71: out <= 32'hA3A3FE5D;
        8'h72: out <= 32'h4040C080;
        8'h73: out <= 32'h8F8F8A05;
        8'h74: out <= 32'h9292AD3F;
        8'h75: out <= 32'h9D9DBC21;
        8'h76: out <= 32'h38384870;
        8'h77: out <= 32'hF5F504F1;
        8'h78: out <= 32'hBCBCDF63;
        8'h79: out <= 32'hB6B6C177;
        8'h7A: out <= 32'hDADA75AF;
        8'h7B: out <= 32'h21216342;
        8'h7C: out <= 32'h10103020;
        8'h7D: out <= 32'hFFFF1AE5;
        8'h7E: out <= 32'hF3F30EFD;
        8'h7F: out <= 32'hD2D26DBF;
        8'h80: out <= 32'hCDCD4C81;
        8'h81: out <= 32'h0C0C1418;
        8'h82: out <= 32'h13133526;
        8'h83: out <= 32'hECEC2FC3;
        8'h84: out <= 32'h5F5FE1BE;
        8'h85: out <= 32'h9797A235;
        8'h86: out <= 32'h4444CC88;
        8'h87: out <= 32'h1717392E;
        8'h88: out <= 32'hC4C45793;
        8'h89: out <= 32'hA7A7F255;
        8'h8A: out <= 32'h7E7E82FC;
        8'h8B: out <= 32'h3D3D477A;
        8'h8C: out <= 32'h6464ACC8;
        8'h8D: out <= 32'h5D5DE7BA;
        8'h8E: out <= 32'h19192B32;
        8'h8F: out <= 32'h737395E6;
        8'h90: out <= 32'h6060A0C0;
        8'h91: out <= 32'h81819819;
        8'h92: out <= 32'h4F4FD19E;
        8'h93: out <= 32'hDCDC7FA3;
        8'h94: out <= 32'h22226644;
        8'h95: out <= 32'h2A2A7E54;
        8'h96: out <= 32'h9090AB3B;
        8'h97: out <= 32'h8888830B;
        8'h98: out <= 32'h4646CA8C;
        8'h99: out <= 32'hEEEE29C7;
        8'h9A: out <= 32'hB8B8D36B;
        8'h9B: out <= 32'h14143C28;
        8'h9C: out <= 32'hDEDE79A7;
        8'h9D: out <= 32'h5E5EE2BC;
        8'h9E: out <= 32'h0B0B1D16;
        8'h9F: out <= 32'hDBDB76AD;
        8'hA0: out <= 32'hE0E03BDB;
        8'hA1: out <= 32'h32325664;
        8'hA2: out <= 32'h3A3A4E74;
        8'hA3: out <= 32'h0A0A1E14;
        8'hA4: out <= 32'h4949DB92;
        8'hA5: out <= 32'h06060A0C;
        8'hA6: out <= 32'h24246C48;
        8'hA7: out <= 32'h5C5CE4B8;
        8'hA8: out <= 32'hC2C25D9F;
        8'hA9: out <= 32'hD3D36EBD;
        8'hAA: out <= 32'hACACEF43;
        8'hAB: out <= 32'h6262A6C4;
        8'hAC: out <= 32'h9191A839;
        8'hAD: out <= 32'h9595A431;
        8'hAE: out <= 32'hE4E437D3;
        8'hAF: out <= 32'h79798BF2;
        8'hB0: out <= 32'hE7E732D5;
        8'hB1: out <= 32'hC8C8438B;
        8'hB2: out <= 32'h3737596E;
        8'hB3: out <= 32'h6D6DB7DA;
        8'hB4: out <= 32'h8D8D8C01;
        8'hB5: out <= 32'hD5D564B1;
        8'hB6: out <= 32'h4E4ED29C;
        8'hB7: out <= 32'hA9A9E049;
        8'hB8: out <= 32'h6C6CB4D8;
        8'hB9: out <= 32'h5656FAAC;
        8'hBA: out <= 32'hF4F407F3;
        8'hBB: out <= 32'hEAEA25CF;
        8'hBC: out <= 32'h6565AFCA;
        8'hBD: out <= 32'h7A7A8EF4;
        8'hBE: out <= 32'hAEAEE947;
        8'hBF: out <= 32'h08081810;
        8'hC0: out <= 32'hBABAD56F;
        8'hC1: out <= 32'h787888F0;
        8'hC2: out <= 32'h25256F4A;
        8'hC3: out <= 32'h2E2E725C;
        8'hC4: out <= 32'h1C1C2438;
        8'hC5: out <= 32'hA6A6F157;
        8'hC6: out <= 32'hB4B4C773;
        8'hC7: out <= 32'hC6C65197;
        8'hC8: out <= 32'hE8E823CB;
        8'hC9: out <= 32'hDDDD7CA1;
        8'hCA: out <= 32'h74749CE8;
        8'hCB: out <= 32'h1F1F213E;
        8'hCC: out <= 32'h4B4BDD96;
        8'hCD: out <= 32'hBDBDDC61;
        8'hCE: out <= 32'h8B8B860D;
        8'hCF: out <= 32'h8A8A850F;
        8'hD0: out <= 32'h707090E0;
        8'hD1: out <= 32'h3E3E427C;
        8'hD2: out <= 32'hB5B5C471;
        8'hD3: out <= 32'h6666AACC;
        8'hD4: out <= 32'h4848D890;
        8'hD5: out <= 32'h03030506;
        8'hD6: out <= 32'hF6F601F7;
        8'hD7: out <= 32'h0E0E121C;
        8'hD8: out <= 32'h6161A3C2;
        8'hD9: out <= 32'h35355F6A;
        8'hDA: out <= 32'h5757F9AE;
        8'hDB: out <= 32'hB9B9D069;
        8'hDC: out <= 32'h86869117;
        8'hDD: out <= 32'hC1C15899;
        8'hDE: out <= 32'h1D1D273A;
        8'hDF: out <= 32'h9E9EB927;
        8'hE0: out <= 32'hE1E138D9;
        8'hE1: out <= 32'hF8F813EB;
        8'hE2: out <= 32'h9898B32B;
        8'hE3: out <= 32'h11113322;
        8'hE4: out <= 32'h6969BBD2;
        8'hE5: out <= 32'hD9D970A9;
        8'hE6: out <= 32'h8E8E8907;
        8'hE7: out <= 32'h9494A733;
        8'hE8: out <= 32'h9B9BB62D;
        8'hE9: out <= 32'h1E1E223C;
        8'hEA: out <= 32'h87879215;
        8'hEB: out <= 32'hE9E920C9;
        8'hEC: out <= 32'hCECE4987;
        8'hED: out <= 32'h5555FFAA;
        8'hEE: out <= 32'h28287850;
        8'hEF: out <= 32'hDFDF7AA5;
        8'hF0: out <= 32'h8C8C8F03;
        8'hF1: out <= 32'hA1A1F859;
        8'hF2: out <= 32'h89898009;
        8'hF3: out <= 32'h0D0D171A;
        8'hF4: out <= 32'hBFBFDA65;
        8'hF5: out <= 32'hE6E631D7;
        8'hF6: out <= 32'h4242C684;
        8'hF7: out <= 32'h6868B8D0;
        8'hF8: out <= 32'h4141C382;
        8'hF9: out <= 32'h9999B029;
        8'hFA: out <= 32'h2D2D775A;
        8'hFB: out <= 32'h0F0F111E;
        8'hFC: out <= 32'hB0B0CB7B;
        8'hFD: out <= 32'h5454FCA8;
        8'hFE: out <= 32'hBBBBD66D;
        8'hFF: out <= 32'h16163A2C;
        endcase
    end
endmodule
